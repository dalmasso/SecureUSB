------------------------------------------------------------------------
-- Engineer:    Dalmasso Loic
-- Create Date: 25/08/2025
-- Module Name: USBVerifierWrapper
-- Description:
--		The USBVerifier Wrapper Module embedds USBVerifier and all components required to perform USB Verification Field Values
--
-- Ports
--		Input 	-	i_sys_clock: System Input Clock
--		Input 	-	i_enable: System Input Enable ('0': Disabled, '1': Enabled)
--		Input 	-	i_descriptor_field: Descriptor Field to verify
--		Input 	-	i_descriptor_field_available: Descriptor Field Available ('0': Not Available, '1': Available)
--		Input 	-	i_descriptor_value: Descriptor Value to verify
--		Input 	-	i_descriptor_value_en: Descriptor Value Quartet Enable ('0': Disabled Quartet, '1': Enabled Quartet)
--		Input 	-	i_descriptor_value_total_part_number: Descriptor Value Total Part Number to verify
--		Input 	-	i_descriptor_value_part_number: Descriptor Value Part Number to verify
--		Input 	-	i_descriptor_value_new_part: New Descriptor Value Part ('0': No New Part, '1': New Part)
--		Output 	-	o_descriptor_value_next_part_request: Next Descriptor Value Part Request ('0': No Request, '1': New Request)
--		Output 	-	o_ready: Verification Result Ready ('0': Not Ready, '1': Ready)
--		Output 	-	o_result: Verification Result ('0': Error, '1': Success)
------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

-- Custom Package: USB Descriptor Fields
LIBRARY WORK;
USE WORK.USBDescriptorFields.ALL;

-- Custom Package: USB Descriptor Values
LIBRARY WORK;
USE WORK.USBDescriptorValues.ALL;

ENTITY USBVerifierWrapper is

PORT(
	i_sys_clock: IN STD_LOGIC;
	i_enable: IN STD_LOGIC;
	i_descriptor_field: IN UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0);
	i_descriptor_field_available: IN STD_LOGIC;
	i_descriptor_value: IN UNSIGNED(USB_DESCRIPTOR_VALUE_DATA_BIT_LENGTH-1 downto 0);
	i_descriptor_value_en: IN STD_LOGIC_VECTOR(USB_DESCRIPTOR_VALUE_QUARTET_EN_BIT_LENGTH-1 downto 0);
    i_descriptor_value_total_part_number: IN UNSIGNED(USB_DESCRIPTOR_VALUE_PART_NUMBER_BIT_LENGTH-1 downto 0);
	i_descriptor_value_part_number: IN UNSIGNED(USB_DESCRIPTOR_VALUE_PART_NUMBER_BIT_LENGTH-1 downto 0);
	i_descriptor_value_new_part: IN STD_LOGIC;
	o_descriptor_value_next_part_request: OUT STD_LOGIC;
	o_ready: OUT STD_LOGIC;
	o_result: OUT STD_LOGIC
);

END USBVerifierWrapper;

ARCHITECTURE Behavioral of USBVerifierWrapper is

------------------------------------------------------------------------
-- Component Declarations
------------------------------------------------------------------------
COMPONENT USBVerifier is
GENERIC(
	EQUALS_OPERATOR_ENABLE: STD_LOGIC := '1';
	NOT_EQUALS_OPERATOR_ENABLE: STD_LOGIC := '1';
	GREATER_OPERATOR_ENABLE: STD_LOGIC := '1';
	GREATER_EQUALS_OPERATOR_ENABLE: STD_LOGIC := '1';
	LESS_OPERATOR_ENABLE: STD_LOGIC := '1';
	LESS_EQUALS_OPERATOR_ENABLE: STD_LOGIC := '1';
	STARTS_WITH_OPERATOR_ENABLE: STD_LOGIC := '1';
	ENDS_WITH_OPERATOR_ENABLE: STD_LOGIC := '1';
	CONTAINS_OPERATOR_ENABLE: STD_LOGIC := '1';
	NOT_CONTAINS_OPERATOR_ENABLE: STD_LOGIC := '1';
	WATCHDOG_LIMIT: INTEGER := 18;

	EQUALS_MEMORY_ADDR_LENGTH: INTEGER := 1;
	EQUALS_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	EQUALS_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	EQUALS_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	EQUALS_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	EQUALS_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	EQUALS_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	EQUALS_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	EQUALS_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	EQUALS_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	EQUALS_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	EQUALS_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	EQUALS_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	EQUALS_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	EQUALS_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	EQUALS_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	EQUALS_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	EQUALS_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	EQUALS_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	EQUALS_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	EQUALS_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	EQUALS_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	EQUALS_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	EQUALS_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	EQUALS_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	EQUALS_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	EQUALS_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	EQUALS_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	EQUALS_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	EQUALS_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	EQUALS_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	EQUALS_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	EQUALS_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	EQUALS_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	EQUALS_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	EQUALS_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	EQUALS_HID_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_HID_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_HID_BCDHID_INDEX: INTEGER := 0;
	EQUALS_HID_BCDHID_COUNT: INTEGER := 0;
	EQUALS_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	EQUALS_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	EQUALS_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	EQUALS_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	EQUALS_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	EQUALS_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	EQUALS_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	EQUALS_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	EQUALS_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	EQUALS_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	EQUALS_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	EQUALS_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	EQUALS_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	EQUALS_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	EQUALS_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	EQUALS_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	EQUALS_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	EQUALS_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	EQUALS_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	EQUALS_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	EQUALS_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	EQUALS_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	EQUALS_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	EQUALS_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	EQUALS_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	EQUALS_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	EQUALS_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	NOT_EQUALS_MEMORY_ADDR_LENGTH: INTEGER := 1;
	NOT_EQUALS_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	NOT_EQUALS_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	NOT_EQUALS_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	NOT_EQUALS_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	NOT_EQUALS_HID_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_HID_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_HID_BCDHID_INDEX: INTEGER := 0;
	NOT_EQUALS_HID_BCDHID_COUNT: INTEGER := 0;
	NOT_EQUALS_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	NOT_EQUALS_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	NOT_EQUALS_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	NOT_EQUALS_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	NOT_EQUALS_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	NOT_EQUALS_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	NOT_EQUALS_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	NOT_EQUALS_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	NOT_EQUALS_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	NOT_EQUALS_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	GREATER_MEMORY_ADDR_LENGTH: INTEGER := 1;
	GREATER_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	GREATER_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	GREATER_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	GREATER_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	GREATER_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	GREATER_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	GREATER_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	GREATER_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	GREATER_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	GREATER_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	GREATER_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	GREATER_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	GREATER_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	GREATER_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	GREATER_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	GREATER_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	GREATER_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	GREATER_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	GREATER_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	GREATER_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	GREATER_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	GREATER_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	GREATER_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	GREATER_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	GREATER_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	GREATER_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	GREATER_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	GREATER_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	GREATER_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	GREATER_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	GREATER_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	GREATER_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	GREATER_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	GREATER_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	GREATER_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	GREATER_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	GREATER_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	GREATER_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	GREATER_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	GREATER_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	GREATER_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	GREATER_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	GREATER_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	GREATER_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	GREATER_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	GREATER_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	GREATER_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	GREATER_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	GREATER_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	GREATER_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	GREATER_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	GREATER_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	GREATER_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	GREATER_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	GREATER_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	GREATER_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	GREATER_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	GREATER_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	GREATER_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	GREATER_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	GREATER_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	GREATER_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	GREATER_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	GREATER_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	GREATER_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	GREATER_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	GREATER_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	GREATER_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	GREATER_HID_BLENGTH_INDEX: INTEGER := 0;
	GREATER_HID_BLENGTH_COUNT: INTEGER := 0;
	GREATER_HID_BCDHID_INDEX: INTEGER := 0;
	GREATER_HID_BCDHID_COUNT: INTEGER := 0;
	GREATER_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	GREATER_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	GREATER_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	GREATER_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	GREATER_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	GREATER_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	GREATER_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	GREATER_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	GREATER_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	GREATER_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	GREATER_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	GREATER_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	GREATER_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	GREATER_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	GREATER_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	GREATER_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	GREATER_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	GREATER_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	GREATER_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	GREATER_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	GREATER_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	GREATER_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	GREATER_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	GREATER_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	GREATER_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	GREATER_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	GREATER_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	GREATER_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	GREATER_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	GREATER_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	GREATER_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	GREATER_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	GREATER_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	GREATER_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	GREATER_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	GREATER_EQUALS_MEMORY_ADDR_LENGTH: INTEGER := 1;
	GREATER_EQUALS_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	GREATER_EQUALS_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	GREATER_EQUALS_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	GREATER_EQUALS_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	GREATER_EQUALS_HID_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_HID_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_HID_BCDHID_INDEX: INTEGER := 0;
	GREATER_EQUALS_HID_BCDHID_COUNT: INTEGER := 0;
	GREATER_EQUALS_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	GREATER_EQUALS_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	GREATER_EQUALS_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	GREATER_EQUALS_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	GREATER_EQUALS_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	GREATER_EQUALS_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	GREATER_EQUALS_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	GREATER_EQUALS_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	GREATER_EQUALS_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	GREATER_EQUALS_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	LESS_MEMORY_ADDR_LENGTH: INTEGER := 1;
	LESS_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	LESS_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	LESS_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	LESS_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	LESS_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	LESS_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	LESS_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	LESS_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	LESS_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	LESS_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	LESS_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	LESS_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	LESS_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	LESS_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	LESS_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	LESS_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	LESS_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	LESS_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	LESS_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	LESS_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	LESS_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	LESS_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	LESS_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	LESS_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	LESS_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	LESS_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	LESS_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	LESS_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	LESS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	LESS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	LESS_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	LESS_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	LESS_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	LESS_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	LESS_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	LESS_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	LESS_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	LESS_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	LESS_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	LESS_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	LESS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	LESS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	LESS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	LESS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	LESS_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	LESS_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	LESS_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	LESS_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	LESS_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	LESS_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	LESS_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	LESS_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	LESS_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	LESS_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	LESS_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	LESS_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	LESS_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	LESS_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	LESS_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	LESS_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	LESS_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	LESS_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	LESS_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	LESS_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	LESS_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	LESS_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	LESS_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	LESS_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	LESS_HID_BLENGTH_INDEX: INTEGER := 0;
	LESS_HID_BLENGTH_COUNT: INTEGER := 0;
	LESS_HID_BCDHID_INDEX: INTEGER := 0;
	LESS_HID_BCDHID_COUNT: INTEGER := 0;
	LESS_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	LESS_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	LESS_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	LESS_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	LESS_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	LESS_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	LESS_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	LESS_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	LESS_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	LESS_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	LESS_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	LESS_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	LESS_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	LESS_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	LESS_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	LESS_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	LESS_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	LESS_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	LESS_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	LESS_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	LESS_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	LESS_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	LESS_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	LESS_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	LESS_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	LESS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	LESS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	LESS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	LESS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	LESS_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	LESS_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	LESS_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	LESS_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	LESS_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	LESS_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	LESS_EQUALS_MEMORY_ADDR_LENGTH: INTEGER := 1;
	LESS_EQUALS_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	LESS_EQUALS_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	LESS_EQUALS_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	LESS_EQUALS_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	LESS_EQUALS_HID_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_HID_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_HID_BCDHID_INDEX: INTEGER := 0;
	LESS_EQUALS_HID_BCDHID_COUNT: INTEGER := 0;
	LESS_EQUALS_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	LESS_EQUALS_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	LESS_EQUALS_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	LESS_EQUALS_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	LESS_EQUALS_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	LESS_EQUALS_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	LESS_EQUALS_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	LESS_EQUALS_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	LESS_EQUALS_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	LESS_EQUALS_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	STARTS_WITH_MEMORY_ADDR_LENGTH: INTEGER := 1;
	STARTS_WITH_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	STARTS_WITH_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	STARTS_WITH_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	STARTS_WITH_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	STARTS_WITH_HID_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_HID_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_HID_BCDHID_INDEX: INTEGER := 0;
	STARTS_WITH_HID_BCDHID_COUNT: INTEGER := 0;
	STARTS_WITH_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	STARTS_WITH_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	STARTS_WITH_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	STARTS_WITH_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	STARTS_WITH_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	STARTS_WITH_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	STARTS_WITH_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	STARTS_WITH_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	STARTS_WITH_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	STARTS_WITH_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	STARTS_WITH_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	STARTS_WITH_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	STARTS_WITH_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	STARTS_WITH_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	STARTS_WITH_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	STARTS_WITH_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	ENDS_WITH_MEMORY_ADDR_LENGTH: INTEGER := 1;
	ENDS_WITH_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	ENDS_WITH_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	ENDS_WITH_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	ENDS_WITH_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	ENDS_WITH_HID_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_HID_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_HID_BCDHID_INDEX: INTEGER := 0;
	ENDS_WITH_HID_BCDHID_COUNT: INTEGER := 0;
	ENDS_WITH_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	ENDS_WITH_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	ENDS_WITH_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	ENDS_WITH_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	ENDS_WITH_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	ENDS_WITH_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	ENDS_WITH_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	ENDS_WITH_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	ENDS_WITH_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	ENDS_WITH_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	ENDS_WITH_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	ENDS_WITH_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	ENDS_WITH_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	ENDS_WITH_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	ENDS_WITH_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	ENDS_WITH_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	CONTAINS_MEMORY_ADDR_LENGTH: INTEGER := 1;
	CONTAINS_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	CONTAINS_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	CONTAINS_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	CONTAINS_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	CONTAINS_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	CONTAINS_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	CONTAINS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	CONTAINS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	CONTAINS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	CONTAINS_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	CONTAINS_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	CONTAINS_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	CONTAINS_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	CONTAINS_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	CONTAINS_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	CONTAINS_HID_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_HID_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_HID_BCDHID_INDEX: INTEGER := 0;
	CONTAINS_HID_BCDHID_COUNT: INTEGER := 0;
	CONTAINS_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	CONTAINS_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	CONTAINS_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	CONTAINS_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	CONTAINS_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	CONTAINS_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	CONTAINS_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	CONTAINS_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	CONTAINS_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	CONTAINS_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	CONTAINS_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	CONTAINS_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	CONTAINS_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	CONTAINS_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	CONTAINS_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	CONTAINS_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	CONTAINS_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	CONTAINS_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	CONTAINS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	CONTAINS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	CONTAINS_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	CONTAINS_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	CONTAINS_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0;

	NOT_CONTAINS_MEMORY_ADDR_LENGTH: INTEGER := 1;
	NOT_CONTAINS_MEMORY_ADDR_MAX_INDEX: INTEGER := 0;
	NOT_CONTAINS_MEMORY_ADDR_MAX_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BCDUSB_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BCDUSB_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BDEVICECLASS_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BDEVICECLASS_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IDVENDOR_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IDVENDOR_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IDPRODUCT_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IDPRODUCT_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BCDDEVICE_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BCDDEVICE_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IMANUFACTURER_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IMANUFACTURER_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IMANUFACTURER_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IMANUFACTURER_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IPRODUCT_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IPRODUCT_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IPRODUCT_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_IPRODUCT_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_ISERIALNUMBER_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_ISERIALNUMBER_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_WTOTALLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_WTOTALLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BNUMINTERFACES_INDEX: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BNUMINTERFACES_COUNT: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_ICONFIGURATION_INDEX: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_ICONFIGURATION_COUNT: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BMATTRIBUTES_INDEX: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BMATTRIBUTES_COUNT: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BMAXPOWER_INDEX: INTEGER := 0;
	NOT_CONTAINS_CONFIGURATION_BMAXPOWER_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BINTERFACENUMBER_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BINTERFACENUMBER_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BALTERNATESETTING_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BALTERNATESETTING_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BNUMENDPOINTS_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BNUMENDPOINTS_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BINTERFACECLASS_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BINTERFACECLASS_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BINTERFACESUBCLASS_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BINTERFACESUBCLASS_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BINTERFACEPROTOCOL_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_BINTERFACEPROTOCOL_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_IINTERFACE_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_IINTERFACE_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_IINTERFACE_INDEX: INTEGER := 0;
	NOT_CONTAINS_INTERFACE_IINTERFACE_COUNT: INTEGER := 0;
	NOT_CONTAINS_HID_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_HID_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_HID_BCDHID_INDEX: INTEGER := 0;
	NOT_CONTAINS_HID_BCDHID_COUNT: INTEGER := 0;
	NOT_CONTAINS_HID_BCOUNTRYCODE_INDEX: INTEGER := 0;
	NOT_CONTAINS_HID_BCOUNTRYCODE_COUNT: INTEGER := 0;
	NOT_CONTAINS_HID_BNUMDESCRIPTORS_INDEX: INTEGER := 0;
	NOT_CONTAINS_HID_BNUMDESCRIPTORS_COUNT: INTEGER := 0;
	NOT_CONTAINS_HID_BDESCRIPTORTYPE_INDEX: INTEGER := 0;
	NOT_CONTAINS_HID_BDESCRIPTORTYPE_COUNT: INTEGER := 0;
	NOT_CONTAINS_HID_WDESCRIPTORLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_HID_WDESCRIPTORLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_BENDPOINTADDRESS_INDEX: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_BENDPOINTADDRESS_COUNT: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_BMATTRIBUTES_INDEX: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_BMATTRIBUTES_COUNT: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_WMAXPACKETSIZE_INDEX: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_WMAXPACKETSIZE_COUNT: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_BINTERVAL_INDEX: INTEGER := 0;
	NOT_CONTAINS_ENDPOINT_BINTERVAL_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BCDUSB_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BCDUSB_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BRESERVED_INDEX: INTEGER := 0;
	NOT_CONTAINS_DEVICE_QUALIFIER_BRESERVED_COUNT: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_WTOTALLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_WTOTALLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BNUMINTERFACES_INDEX: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BNUMINTERFACES_COUNT: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_ICONFIGURATION_INDEX: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_ICONFIGURATION_COUNT: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BMATTRIBUTES_INDEX: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BMATTRIBUTES_COUNT: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BMAXPOWER_INDEX: INTEGER := 0;
	NOT_CONTAINS_OTHER_SPEED_BMAXPOWER_COUNT: INTEGER := 0
);

PORT(
	i_sys_clock: IN STD_LOGIC;
	i_enable: IN STD_LOGIC;
	i_descriptor_field: IN UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0);
	i_descriptor_field_available: IN STD_LOGIC;
	i_descriptor_value: IN UNSIGNED(USB_DESCRIPTOR_VALUE_DATA_BIT_LENGTH-1 downto 0);
	i_descriptor_value_en: IN STD_LOGIC_VECTOR(USB_DESCRIPTOR_VALUE_QUARTET_EN_BIT_LENGTH-1 downto 0);
    i_descriptor_value_total_part_number: IN UNSIGNED(USB_DESCRIPTOR_VALUE_PART_NUMBER_BIT_LENGTH-1 downto 0);
	i_descriptor_value_part_number: IN UNSIGNED(USB_DESCRIPTOR_VALUE_PART_NUMBER_BIT_LENGTH-1 downto 0);
	i_descriptor_value_new_part: IN STD_LOGIC;
	o_descriptor_value_next_part_request: OUT STD_LOGIC;
	o_ready: OUT STD_LOGIC;
	o_result: OUT STD_LOGIC
);

END COMPONENT;

------------------------------------------------------------------------
-- Module Implementation
------------------------------------------------------------------------
begin

	------------------
	-- USB Verifier --
	------------------
	usbVerifier_inst: USBVerifier
		GENERIC MAP (
			EQUALS_OPERATOR_ENABLE => '1',
			NOT_EQUALS_OPERATOR_ENABLE => '1',
			GREATER_OPERATOR_ENABLE => '1',
			GREATER_EQUALS_OPERATOR_ENABLE => '1',
			LESS_OPERATOR_ENABLE => '1',
			LESS_EQUALS_OPERATOR_ENABLE => '1',
			STARTS_WITH_OPERATOR_ENABLE => '1',
			ENDS_WITH_OPERATOR_ENABLE => '1',
			CONTAINS_OPERATOR_ENABLE => '1',
			NOT_CONTAINS_OPERATOR_ENABLE => '1',
			WATCHDOG_LIMIT => 18,

			EQUALS_MEMORY_ADDR_LENGTH => 1,
			EQUALS_MEMORY_ADDR_MAX_INDEX => 0,
			EQUALS_MEMORY_ADDR_MAX_COUNT => 0,
			EQUALS_DEVICE_BLENGTH_INDEX => 0,
			EQUALS_DEVICE_BLENGTH_COUNT => 0,
			EQUALS_DEVICE_BCDUSB_INDEX => 0,
			EQUALS_DEVICE_BCDUSB_COUNT => 0,
			EQUALS_DEVICE_BDEVICECLASS_INDEX => 0,
			EQUALS_DEVICE_BDEVICECLASS_COUNT => 0,
			EQUALS_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			EQUALS_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			EQUALS_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			EQUALS_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			EQUALS_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			EQUALS_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			EQUALS_DEVICE_IDVENDOR_INDEX => 0,
			EQUALS_DEVICE_IDVENDOR_COUNT => 0,
			EQUALS_DEVICE_IDPRODUCT_INDEX => 0,
			EQUALS_DEVICE_IDPRODUCT_COUNT => 0,
			EQUALS_DEVICE_BCDDEVICE_INDEX => 0,
			EQUALS_DEVICE_BCDDEVICE_COUNT => 0,
			EQUALS_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			EQUALS_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			EQUALS_DEVICE_IMANUFACTURER_INDEX => 0,
			EQUALS_DEVICE_IMANUFACTURER_COUNT => 0,
			EQUALS_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			EQUALS_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			EQUALS_DEVICE_IPRODUCT_INDEX => 0,
			EQUALS_DEVICE_IPRODUCT_COUNT => 0,
			EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			EQUALS_DEVICE_ISERIALNUMBER_INDEX => 0,
			EQUALS_DEVICE_ISERIALNUMBER_COUNT => 0,
			EQUALS_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			EQUALS_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			EQUALS_CONFIGURATION_BLENGTH_INDEX => 0,
			EQUALS_CONFIGURATION_BLENGTH_COUNT => 0,
			EQUALS_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			EQUALS_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			EQUALS_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			EQUALS_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			EQUALS_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			EQUALS_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			EQUALS_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			EQUALS_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			EQUALS_CONFIGURATION_BMAXPOWER_INDEX => 0,
			EQUALS_CONFIGURATION_BMAXPOWER_COUNT => 0,
			EQUALS_INTERFACE_BLENGTH_INDEX => 0,
			EQUALS_INTERFACE_BLENGTH_COUNT => 0,
			EQUALS_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			EQUALS_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			EQUALS_INTERFACE_BALTERNATESETTING_INDEX => 0,
			EQUALS_INTERFACE_BALTERNATESETTING_COUNT => 0,
			EQUALS_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			EQUALS_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			EQUALS_INTERFACE_BINTERFACECLASS_INDEX => 0,
			EQUALS_INTERFACE_BINTERFACECLASS_COUNT => 0,
			EQUALS_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			EQUALS_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			EQUALS_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			EQUALS_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			EQUALS_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			EQUALS_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			EQUALS_INTERFACE_IINTERFACE_INDEX => 0,
			EQUALS_INTERFACE_IINTERFACE_COUNT => 0,
			EQUALS_HID_BLENGTH_INDEX => 0,
			EQUALS_HID_BLENGTH_COUNT => 0,
			EQUALS_HID_BCDHID_INDEX => 0,
			EQUALS_HID_BCDHID_COUNT => 0,
			EQUALS_HID_BCOUNTRYCODE_INDEX => 0,
			EQUALS_HID_BCOUNTRYCODE_COUNT => 0,
			EQUALS_HID_BNUMDESCRIPTORS_INDEX => 0,
			EQUALS_HID_BNUMDESCRIPTORS_COUNT => 0,
			EQUALS_HID_BDESCRIPTORTYPE_INDEX => 0,
			EQUALS_HID_BDESCRIPTORTYPE_COUNT => 0,
			EQUALS_HID_WDESCRIPTORLENGTH_INDEX => 0,
			EQUALS_HID_WDESCRIPTORLENGTH_COUNT => 0,
			EQUALS_ENDPOINT_BLENGTH_INDEX => 0,
			EQUALS_ENDPOINT_BLENGTH_COUNT => 0,
			EQUALS_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			EQUALS_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			EQUALS_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			EQUALS_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			EQUALS_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			EQUALS_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			EQUALS_ENDPOINT_BINTERVAL_INDEX => 0,
			EQUALS_ENDPOINT_BINTERVAL_COUNT => 0,
			EQUALS_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			EQUALS_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			EQUALS_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			EQUALS_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			EQUALS_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			EQUALS_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			EQUALS_OTHER_SPEED_BLENGTH_INDEX => 0,
			EQUALS_OTHER_SPEED_BLENGTH_COUNT => 0,
			EQUALS_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			EQUALS_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			EQUALS_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			EQUALS_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			EQUALS_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			EQUALS_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			EQUALS_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			EQUALS_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			EQUALS_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			EQUALS_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			NOT_EQUALS_MEMORY_ADDR_LENGTH => 1,
			NOT_EQUALS_MEMORY_ADDR_MAX_INDEX => 0,
			NOT_EQUALS_MEMORY_ADDR_MAX_COUNT => 0,
			NOT_EQUALS_DEVICE_BLENGTH_INDEX => 0,
			NOT_EQUALS_DEVICE_BLENGTH_COUNT => 0,
			NOT_EQUALS_DEVICE_BCDUSB_INDEX => 0,
			NOT_EQUALS_DEVICE_BCDUSB_COUNT => 0,
			NOT_EQUALS_DEVICE_BDEVICECLASS_INDEX => 0,
			NOT_EQUALS_DEVICE_BDEVICECLASS_COUNT => 0,
			NOT_EQUALS_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			NOT_EQUALS_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			NOT_EQUALS_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			NOT_EQUALS_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			NOT_EQUALS_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			NOT_EQUALS_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			NOT_EQUALS_DEVICE_IDVENDOR_INDEX => 0,
			NOT_EQUALS_DEVICE_IDVENDOR_COUNT => 0,
			NOT_EQUALS_DEVICE_IDPRODUCT_INDEX => 0,
			NOT_EQUALS_DEVICE_IDPRODUCT_COUNT => 0,
			NOT_EQUALS_DEVICE_BCDDEVICE_INDEX => 0,
			NOT_EQUALS_DEVICE_BCDDEVICE_COUNT => 0,
			NOT_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			NOT_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			NOT_EQUALS_DEVICE_IMANUFACTURER_INDEX => 0,
			NOT_EQUALS_DEVICE_IMANUFACTURER_COUNT => 0,
			NOT_EQUALS_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			NOT_EQUALS_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			NOT_EQUALS_DEVICE_IPRODUCT_INDEX => 0,
			NOT_EQUALS_DEVICE_IPRODUCT_COUNT => 0,
			NOT_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			NOT_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			NOT_EQUALS_DEVICE_ISERIALNUMBER_INDEX => 0,
			NOT_EQUALS_DEVICE_ISERIALNUMBER_COUNT => 0,
			NOT_EQUALS_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			NOT_EQUALS_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			NOT_EQUALS_CONFIGURATION_BLENGTH_INDEX => 0,
			NOT_EQUALS_CONFIGURATION_BLENGTH_COUNT => 0,
			NOT_EQUALS_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			NOT_EQUALS_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			NOT_EQUALS_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			NOT_EQUALS_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			NOT_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			NOT_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			NOT_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			NOT_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			NOT_EQUALS_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			NOT_EQUALS_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			NOT_EQUALS_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			NOT_EQUALS_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			NOT_EQUALS_CONFIGURATION_BMAXPOWER_INDEX => 0,
			NOT_EQUALS_CONFIGURATION_BMAXPOWER_COUNT => 0,
			NOT_EQUALS_INTERFACE_BLENGTH_INDEX => 0,
			NOT_EQUALS_INTERFACE_BLENGTH_COUNT => 0,
			NOT_EQUALS_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			NOT_EQUALS_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			NOT_EQUALS_INTERFACE_BALTERNATESETTING_INDEX => 0,
			NOT_EQUALS_INTERFACE_BALTERNATESETTING_COUNT => 0,
			NOT_EQUALS_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			NOT_EQUALS_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			NOT_EQUALS_INTERFACE_BINTERFACECLASS_INDEX => 0,
			NOT_EQUALS_INTERFACE_BINTERFACECLASS_COUNT => 0,
			NOT_EQUALS_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			NOT_EQUALS_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			NOT_EQUALS_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			NOT_EQUALS_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			NOT_EQUALS_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			NOT_EQUALS_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			NOT_EQUALS_INTERFACE_IINTERFACE_INDEX => 0,
			NOT_EQUALS_INTERFACE_IINTERFACE_COUNT => 0,
			NOT_EQUALS_HID_BLENGTH_INDEX => 0,
			NOT_EQUALS_HID_BLENGTH_COUNT => 0,
			NOT_EQUALS_HID_BCDHID_INDEX => 0,
			NOT_EQUALS_HID_BCDHID_COUNT => 0,
			NOT_EQUALS_HID_BCOUNTRYCODE_INDEX => 0,
			NOT_EQUALS_HID_BCOUNTRYCODE_COUNT => 0,
			NOT_EQUALS_HID_BNUMDESCRIPTORS_INDEX => 0,
			NOT_EQUALS_HID_BNUMDESCRIPTORS_COUNT => 0,
			NOT_EQUALS_HID_BDESCRIPTORTYPE_INDEX => 0,
			NOT_EQUALS_HID_BDESCRIPTORTYPE_COUNT => 0,
			NOT_EQUALS_HID_WDESCRIPTORLENGTH_INDEX => 0,
			NOT_EQUALS_HID_WDESCRIPTORLENGTH_COUNT => 0,
			NOT_EQUALS_ENDPOINT_BLENGTH_INDEX => 0,
			NOT_EQUALS_ENDPOINT_BLENGTH_COUNT => 0,
			NOT_EQUALS_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			NOT_EQUALS_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			NOT_EQUALS_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			NOT_EQUALS_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			NOT_EQUALS_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			NOT_EQUALS_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			NOT_EQUALS_ENDPOINT_BINTERVAL_INDEX => 0,
			NOT_EQUALS_ENDPOINT_BINTERVAL_COUNT => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			NOT_EQUALS_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			NOT_EQUALS_OTHER_SPEED_BLENGTH_INDEX => 0,
			NOT_EQUALS_OTHER_SPEED_BLENGTH_COUNT => 0,
			NOT_EQUALS_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			NOT_EQUALS_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			NOT_EQUALS_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			NOT_EQUALS_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			NOT_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			NOT_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			NOT_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			NOT_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			NOT_EQUALS_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			NOT_EQUALS_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			NOT_EQUALS_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			NOT_EQUALS_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			NOT_EQUALS_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			NOT_EQUALS_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			GREATER_MEMORY_ADDR_LENGTH => 1,
			GREATER_MEMORY_ADDR_MAX_INDEX => 0,
			GREATER_MEMORY_ADDR_MAX_COUNT => 0,
			GREATER_DEVICE_BLENGTH_INDEX => 0,
			GREATER_DEVICE_BLENGTH_COUNT => 0,
			GREATER_DEVICE_BCDUSB_INDEX => 0,
			GREATER_DEVICE_BCDUSB_COUNT => 0,
			GREATER_DEVICE_BDEVICECLASS_INDEX => 0,
			GREATER_DEVICE_BDEVICECLASS_COUNT => 0,
			GREATER_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			GREATER_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			GREATER_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			GREATER_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			GREATER_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			GREATER_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			GREATER_DEVICE_IDVENDOR_INDEX => 0,
			GREATER_DEVICE_IDVENDOR_COUNT => 0,
			GREATER_DEVICE_IDPRODUCT_INDEX => 0,
			GREATER_DEVICE_IDPRODUCT_COUNT => 0,
			GREATER_DEVICE_BCDDEVICE_INDEX => 0,
			GREATER_DEVICE_BCDDEVICE_COUNT => 0,
			GREATER_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			GREATER_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			GREATER_DEVICE_IMANUFACTURER_INDEX => 0,
			GREATER_DEVICE_IMANUFACTURER_COUNT => 0,
			GREATER_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			GREATER_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			GREATER_DEVICE_IPRODUCT_INDEX => 0,
			GREATER_DEVICE_IPRODUCT_COUNT => 0,
			GREATER_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			GREATER_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			GREATER_DEVICE_ISERIALNUMBER_INDEX => 0,
			GREATER_DEVICE_ISERIALNUMBER_COUNT => 0,
			GREATER_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			GREATER_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			GREATER_CONFIGURATION_BLENGTH_INDEX => 0,
			GREATER_CONFIGURATION_BLENGTH_COUNT => 0,
			GREATER_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			GREATER_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			GREATER_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			GREATER_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			GREATER_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			GREATER_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			GREATER_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			GREATER_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			GREATER_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			GREATER_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			GREATER_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			GREATER_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			GREATER_CONFIGURATION_BMAXPOWER_INDEX => 0,
			GREATER_CONFIGURATION_BMAXPOWER_COUNT => 0,
			GREATER_INTERFACE_BLENGTH_INDEX => 0,
			GREATER_INTERFACE_BLENGTH_COUNT => 0,
			GREATER_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			GREATER_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			GREATER_INTERFACE_BALTERNATESETTING_INDEX => 0,
			GREATER_INTERFACE_BALTERNATESETTING_COUNT => 0,
			GREATER_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			GREATER_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			GREATER_INTERFACE_BINTERFACECLASS_INDEX => 0,
			GREATER_INTERFACE_BINTERFACECLASS_COUNT => 0,
			GREATER_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			GREATER_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			GREATER_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			GREATER_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			GREATER_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			GREATER_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			GREATER_INTERFACE_IINTERFACE_INDEX => 0,
			GREATER_INTERFACE_IINTERFACE_COUNT => 0,
			GREATER_HID_BLENGTH_INDEX => 0,
			GREATER_HID_BLENGTH_COUNT => 0,
			GREATER_HID_BCDHID_INDEX => 0,
			GREATER_HID_BCDHID_COUNT => 0,
			GREATER_HID_BCOUNTRYCODE_INDEX => 0,
			GREATER_HID_BCOUNTRYCODE_COUNT => 0,
			GREATER_HID_BNUMDESCRIPTORS_INDEX => 0,
			GREATER_HID_BNUMDESCRIPTORS_COUNT => 0,
			GREATER_HID_BDESCRIPTORTYPE_INDEX => 0,
			GREATER_HID_BDESCRIPTORTYPE_COUNT => 0,
			GREATER_HID_WDESCRIPTORLENGTH_INDEX => 0,
			GREATER_HID_WDESCRIPTORLENGTH_COUNT => 0,
			GREATER_ENDPOINT_BLENGTH_INDEX => 0,
			GREATER_ENDPOINT_BLENGTH_COUNT => 0,
			GREATER_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			GREATER_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			GREATER_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			GREATER_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			GREATER_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			GREATER_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			GREATER_ENDPOINT_BINTERVAL_INDEX => 0,
			GREATER_ENDPOINT_BINTERVAL_COUNT => 0,
			GREATER_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			GREATER_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			GREATER_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			GREATER_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			GREATER_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			GREATER_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			GREATER_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			GREATER_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			GREATER_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			GREATER_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			GREATER_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			GREATER_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			GREATER_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			GREATER_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			GREATER_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			GREATER_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			GREATER_OTHER_SPEED_BLENGTH_INDEX => 0,
			GREATER_OTHER_SPEED_BLENGTH_COUNT => 0,
			GREATER_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			GREATER_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			GREATER_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			GREATER_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			GREATER_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			GREATER_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			GREATER_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			GREATER_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			GREATER_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			GREATER_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			GREATER_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			GREATER_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			GREATER_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			GREATER_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			GREATER_EQUALS_MEMORY_ADDR_LENGTH => 1,
			GREATER_EQUALS_MEMORY_ADDR_MAX_INDEX => 0,
			GREATER_EQUALS_MEMORY_ADDR_MAX_COUNT => 0,
			GREATER_EQUALS_DEVICE_BLENGTH_INDEX => 0,
			GREATER_EQUALS_DEVICE_BLENGTH_COUNT => 0,
			GREATER_EQUALS_DEVICE_BCDUSB_INDEX => 0,
			GREATER_EQUALS_DEVICE_BCDUSB_COUNT => 0,
			GREATER_EQUALS_DEVICE_BDEVICECLASS_INDEX => 0,
			GREATER_EQUALS_DEVICE_BDEVICECLASS_COUNT => 0,
			GREATER_EQUALS_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			GREATER_EQUALS_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			GREATER_EQUALS_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			GREATER_EQUALS_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			GREATER_EQUALS_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			GREATER_EQUALS_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			GREATER_EQUALS_DEVICE_IDVENDOR_INDEX => 0,
			GREATER_EQUALS_DEVICE_IDVENDOR_COUNT => 0,
			GREATER_EQUALS_DEVICE_IDPRODUCT_INDEX => 0,
			GREATER_EQUALS_DEVICE_IDPRODUCT_COUNT => 0,
			GREATER_EQUALS_DEVICE_BCDDEVICE_INDEX => 0,
			GREATER_EQUALS_DEVICE_BCDDEVICE_COUNT => 0,
			GREATER_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			GREATER_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			GREATER_EQUALS_DEVICE_IMANUFACTURER_INDEX => 0,
			GREATER_EQUALS_DEVICE_IMANUFACTURER_COUNT => 0,
			GREATER_EQUALS_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			GREATER_EQUALS_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			GREATER_EQUALS_DEVICE_IPRODUCT_INDEX => 0,
			GREATER_EQUALS_DEVICE_IPRODUCT_COUNT => 0,
			GREATER_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			GREATER_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			GREATER_EQUALS_DEVICE_ISERIALNUMBER_INDEX => 0,
			GREATER_EQUALS_DEVICE_ISERIALNUMBER_COUNT => 0,
			GREATER_EQUALS_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			GREATER_EQUALS_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			GREATER_EQUALS_CONFIGURATION_BLENGTH_INDEX => 0,
			GREATER_EQUALS_CONFIGURATION_BLENGTH_COUNT => 0,
			GREATER_EQUALS_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			GREATER_EQUALS_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			GREATER_EQUALS_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			GREATER_EQUALS_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			GREATER_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			GREATER_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			GREATER_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			GREATER_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			GREATER_EQUALS_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			GREATER_EQUALS_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			GREATER_EQUALS_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			GREATER_EQUALS_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			GREATER_EQUALS_CONFIGURATION_BMAXPOWER_INDEX => 0,
			GREATER_EQUALS_CONFIGURATION_BMAXPOWER_COUNT => 0,
			GREATER_EQUALS_INTERFACE_BLENGTH_INDEX => 0,
			GREATER_EQUALS_INTERFACE_BLENGTH_COUNT => 0,
			GREATER_EQUALS_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			GREATER_EQUALS_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			GREATER_EQUALS_INTERFACE_BALTERNATESETTING_INDEX => 0,
			GREATER_EQUALS_INTERFACE_BALTERNATESETTING_COUNT => 0,
			GREATER_EQUALS_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			GREATER_EQUALS_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			GREATER_EQUALS_INTERFACE_BINTERFACECLASS_INDEX => 0,
			GREATER_EQUALS_INTERFACE_BINTERFACECLASS_COUNT => 0,
			GREATER_EQUALS_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			GREATER_EQUALS_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			GREATER_EQUALS_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			GREATER_EQUALS_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			GREATER_EQUALS_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			GREATER_EQUALS_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			GREATER_EQUALS_INTERFACE_IINTERFACE_INDEX => 0,
			GREATER_EQUALS_INTERFACE_IINTERFACE_COUNT => 0,
			GREATER_EQUALS_HID_BLENGTH_INDEX => 0,
			GREATER_EQUALS_HID_BLENGTH_COUNT => 0,
			GREATER_EQUALS_HID_BCDHID_INDEX => 0,
			GREATER_EQUALS_HID_BCDHID_COUNT => 0,
			GREATER_EQUALS_HID_BCOUNTRYCODE_INDEX => 0,
			GREATER_EQUALS_HID_BCOUNTRYCODE_COUNT => 0,
			GREATER_EQUALS_HID_BNUMDESCRIPTORS_INDEX => 0,
			GREATER_EQUALS_HID_BNUMDESCRIPTORS_COUNT => 0,
			GREATER_EQUALS_HID_BDESCRIPTORTYPE_INDEX => 0,
			GREATER_EQUALS_HID_BDESCRIPTORTYPE_COUNT => 0,
			GREATER_EQUALS_HID_WDESCRIPTORLENGTH_INDEX => 0,
			GREATER_EQUALS_HID_WDESCRIPTORLENGTH_COUNT => 0,
			GREATER_EQUALS_ENDPOINT_BLENGTH_INDEX => 0,
			GREATER_EQUALS_ENDPOINT_BLENGTH_COUNT => 0,
			GREATER_EQUALS_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			GREATER_EQUALS_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			GREATER_EQUALS_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			GREATER_EQUALS_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			GREATER_EQUALS_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			GREATER_EQUALS_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			GREATER_EQUALS_ENDPOINT_BINTERVAL_INDEX => 0,
			GREATER_EQUALS_ENDPOINT_BINTERVAL_COUNT => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			GREATER_EQUALS_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			GREATER_EQUALS_OTHER_SPEED_BLENGTH_INDEX => 0,
			GREATER_EQUALS_OTHER_SPEED_BLENGTH_COUNT => 0,
			GREATER_EQUALS_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			GREATER_EQUALS_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			GREATER_EQUALS_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			GREATER_EQUALS_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			GREATER_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			GREATER_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			GREATER_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			GREATER_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			GREATER_EQUALS_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			GREATER_EQUALS_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			GREATER_EQUALS_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			GREATER_EQUALS_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			GREATER_EQUALS_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			GREATER_EQUALS_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			LESS_MEMORY_ADDR_LENGTH => 1,
			LESS_MEMORY_ADDR_MAX_INDEX => 0,
			LESS_MEMORY_ADDR_MAX_COUNT => 0,
			LESS_DEVICE_BLENGTH_INDEX => 0,
			LESS_DEVICE_BLENGTH_COUNT => 0,
			LESS_DEVICE_BCDUSB_INDEX => 0,
			LESS_DEVICE_BCDUSB_COUNT => 0,
			LESS_DEVICE_BDEVICECLASS_INDEX => 0,
			LESS_DEVICE_BDEVICECLASS_COUNT => 0,
			LESS_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			LESS_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			LESS_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			LESS_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			LESS_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			LESS_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			LESS_DEVICE_IDVENDOR_INDEX => 0,
			LESS_DEVICE_IDVENDOR_COUNT => 0,
			LESS_DEVICE_IDPRODUCT_INDEX => 0,
			LESS_DEVICE_IDPRODUCT_COUNT => 0,
			LESS_DEVICE_BCDDEVICE_INDEX => 0,
			LESS_DEVICE_BCDDEVICE_COUNT => 0,
			LESS_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			LESS_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			LESS_DEVICE_IMANUFACTURER_INDEX => 0,
			LESS_DEVICE_IMANUFACTURER_COUNT => 0,
			LESS_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			LESS_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			LESS_DEVICE_IPRODUCT_INDEX => 0,
			LESS_DEVICE_IPRODUCT_COUNT => 0,
			LESS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			LESS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			LESS_DEVICE_ISERIALNUMBER_INDEX => 0,
			LESS_DEVICE_ISERIALNUMBER_COUNT => 0,
			LESS_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			LESS_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			LESS_CONFIGURATION_BLENGTH_INDEX => 0,
			LESS_CONFIGURATION_BLENGTH_COUNT => 0,
			LESS_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			LESS_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			LESS_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			LESS_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			LESS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			LESS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			LESS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			LESS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			LESS_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			LESS_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			LESS_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			LESS_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			LESS_CONFIGURATION_BMAXPOWER_INDEX => 0,
			LESS_CONFIGURATION_BMAXPOWER_COUNT => 0,
			LESS_INTERFACE_BLENGTH_INDEX => 0,
			LESS_INTERFACE_BLENGTH_COUNT => 0,
			LESS_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			LESS_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			LESS_INTERFACE_BALTERNATESETTING_INDEX => 0,
			LESS_INTERFACE_BALTERNATESETTING_COUNT => 0,
			LESS_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			LESS_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			LESS_INTERFACE_BINTERFACECLASS_INDEX => 0,
			LESS_INTERFACE_BINTERFACECLASS_COUNT => 0,
			LESS_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			LESS_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			LESS_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			LESS_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			LESS_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			LESS_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			LESS_INTERFACE_IINTERFACE_INDEX => 0,
			LESS_INTERFACE_IINTERFACE_COUNT => 0,
			LESS_HID_BLENGTH_INDEX => 0,
			LESS_HID_BLENGTH_COUNT => 0,
			LESS_HID_BCDHID_INDEX => 0,
			LESS_HID_BCDHID_COUNT => 0,
			LESS_HID_BCOUNTRYCODE_INDEX => 0,
			LESS_HID_BCOUNTRYCODE_COUNT => 0,
			LESS_HID_BNUMDESCRIPTORS_INDEX => 0,
			LESS_HID_BNUMDESCRIPTORS_COUNT => 0,
			LESS_HID_BDESCRIPTORTYPE_INDEX => 0,
			LESS_HID_BDESCRIPTORTYPE_COUNT => 0,
			LESS_HID_WDESCRIPTORLENGTH_INDEX => 0,
			LESS_HID_WDESCRIPTORLENGTH_COUNT => 0,
			LESS_ENDPOINT_BLENGTH_INDEX => 0,
			LESS_ENDPOINT_BLENGTH_COUNT => 0,
			LESS_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			LESS_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			LESS_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			LESS_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			LESS_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			LESS_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			LESS_ENDPOINT_BINTERVAL_INDEX => 0,
			LESS_ENDPOINT_BINTERVAL_COUNT => 0,
			LESS_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			LESS_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			LESS_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			LESS_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			LESS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			LESS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			LESS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			LESS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			LESS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			LESS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			LESS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			LESS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			LESS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			LESS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			LESS_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			LESS_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			LESS_OTHER_SPEED_BLENGTH_INDEX => 0,
			LESS_OTHER_SPEED_BLENGTH_COUNT => 0,
			LESS_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			LESS_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			LESS_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			LESS_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			LESS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			LESS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			LESS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			LESS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			LESS_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			LESS_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			LESS_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			LESS_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			LESS_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			LESS_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			LESS_EQUALS_MEMORY_ADDR_LENGTH => 1,
			LESS_EQUALS_MEMORY_ADDR_MAX_INDEX => 0,
			LESS_EQUALS_MEMORY_ADDR_MAX_COUNT => 0,
			LESS_EQUALS_DEVICE_BLENGTH_INDEX => 0,
			LESS_EQUALS_DEVICE_BLENGTH_COUNT => 0,
			LESS_EQUALS_DEVICE_BCDUSB_INDEX => 0,
			LESS_EQUALS_DEVICE_BCDUSB_COUNT => 0,
			LESS_EQUALS_DEVICE_BDEVICECLASS_INDEX => 0,
			LESS_EQUALS_DEVICE_BDEVICECLASS_COUNT => 0,
			LESS_EQUALS_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			LESS_EQUALS_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			LESS_EQUALS_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			LESS_EQUALS_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			LESS_EQUALS_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			LESS_EQUALS_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			LESS_EQUALS_DEVICE_IDVENDOR_INDEX => 0,
			LESS_EQUALS_DEVICE_IDVENDOR_COUNT => 0,
			LESS_EQUALS_DEVICE_IDPRODUCT_INDEX => 0,
			LESS_EQUALS_DEVICE_IDPRODUCT_COUNT => 0,
			LESS_EQUALS_DEVICE_BCDDEVICE_INDEX => 0,
			LESS_EQUALS_DEVICE_BCDDEVICE_COUNT => 0,
			LESS_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			LESS_EQUALS_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			LESS_EQUALS_DEVICE_IMANUFACTURER_INDEX => 0,
			LESS_EQUALS_DEVICE_IMANUFACTURER_COUNT => 0,
			LESS_EQUALS_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			LESS_EQUALS_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			LESS_EQUALS_DEVICE_IPRODUCT_INDEX => 0,
			LESS_EQUALS_DEVICE_IPRODUCT_COUNT => 0,
			LESS_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			LESS_EQUALS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			LESS_EQUALS_DEVICE_ISERIALNUMBER_INDEX => 0,
			LESS_EQUALS_DEVICE_ISERIALNUMBER_COUNT => 0,
			LESS_EQUALS_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			LESS_EQUALS_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			LESS_EQUALS_CONFIGURATION_BLENGTH_INDEX => 0,
			LESS_EQUALS_CONFIGURATION_BLENGTH_COUNT => 0,
			LESS_EQUALS_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			LESS_EQUALS_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			LESS_EQUALS_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			LESS_EQUALS_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			LESS_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			LESS_EQUALS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			LESS_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			LESS_EQUALS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			LESS_EQUALS_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			LESS_EQUALS_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			LESS_EQUALS_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			LESS_EQUALS_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			LESS_EQUALS_CONFIGURATION_BMAXPOWER_INDEX => 0,
			LESS_EQUALS_CONFIGURATION_BMAXPOWER_COUNT => 0,
			LESS_EQUALS_INTERFACE_BLENGTH_INDEX => 0,
			LESS_EQUALS_INTERFACE_BLENGTH_COUNT => 0,
			LESS_EQUALS_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			LESS_EQUALS_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			LESS_EQUALS_INTERFACE_BALTERNATESETTING_INDEX => 0,
			LESS_EQUALS_INTERFACE_BALTERNATESETTING_COUNT => 0,
			LESS_EQUALS_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			LESS_EQUALS_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			LESS_EQUALS_INTERFACE_BINTERFACECLASS_INDEX => 0,
			LESS_EQUALS_INTERFACE_BINTERFACECLASS_COUNT => 0,
			LESS_EQUALS_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			LESS_EQUALS_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			LESS_EQUALS_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			LESS_EQUALS_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			LESS_EQUALS_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			LESS_EQUALS_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			LESS_EQUALS_INTERFACE_IINTERFACE_INDEX => 0,
			LESS_EQUALS_INTERFACE_IINTERFACE_COUNT => 0,
			LESS_EQUALS_HID_BLENGTH_INDEX => 0,
			LESS_EQUALS_HID_BLENGTH_COUNT => 0,
			LESS_EQUALS_HID_BCDHID_INDEX => 0,
			LESS_EQUALS_HID_BCDHID_COUNT => 0,
			LESS_EQUALS_HID_BCOUNTRYCODE_INDEX => 0,
			LESS_EQUALS_HID_BCOUNTRYCODE_COUNT => 0,
			LESS_EQUALS_HID_BNUMDESCRIPTORS_INDEX => 0,
			LESS_EQUALS_HID_BNUMDESCRIPTORS_COUNT => 0,
			LESS_EQUALS_HID_BDESCRIPTORTYPE_INDEX => 0,
			LESS_EQUALS_HID_BDESCRIPTORTYPE_COUNT => 0,
			LESS_EQUALS_HID_WDESCRIPTORLENGTH_INDEX => 0,
			LESS_EQUALS_HID_WDESCRIPTORLENGTH_COUNT => 0,
			LESS_EQUALS_ENDPOINT_BLENGTH_INDEX => 0,
			LESS_EQUALS_ENDPOINT_BLENGTH_COUNT => 0,
			LESS_EQUALS_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			LESS_EQUALS_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			LESS_EQUALS_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			LESS_EQUALS_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			LESS_EQUALS_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			LESS_EQUALS_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			LESS_EQUALS_ENDPOINT_BINTERVAL_INDEX => 0,
			LESS_EQUALS_ENDPOINT_BINTERVAL_COUNT => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			LESS_EQUALS_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			LESS_EQUALS_OTHER_SPEED_BLENGTH_INDEX => 0,
			LESS_EQUALS_OTHER_SPEED_BLENGTH_COUNT => 0,
			LESS_EQUALS_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			LESS_EQUALS_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			LESS_EQUALS_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			LESS_EQUALS_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			LESS_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			LESS_EQUALS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			LESS_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			LESS_EQUALS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			LESS_EQUALS_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			LESS_EQUALS_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			LESS_EQUALS_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			LESS_EQUALS_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			LESS_EQUALS_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			LESS_EQUALS_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			STARTS_WITH_MEMORY_ADDR_LENGTH => 1,
			STARTS_WITH_MEMORY_ADDR_MAX_INDEX => 0,
			STARTS_WITH_MEMORY_ADDR_MAX_COUNT => 0,
			STARTS_WITH_DEVICE_BLENGTH_INDEX => 0,
			STARTS_WITH_DEVICE_BLENGTH_COUNT => 0,
			STARTS_WITH_DEVICE_BCDUSB_INDEX => 0,
			STARTS_WITH_DEVICE_BCDUSB_COUNT => 0,
			STARTS_WITH_DEVICE_BDEVICECLASS_INDEX => 0,
			STARTS_WITH_DEVICE_BDEVICECLASS_COUNT => 0,
			STARTS_WITH_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			STARTS_WITH_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			STARTS_WITH_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			STARTS_WITH_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			STARTS_WITH_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			STARTS_WITH_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			STARTS_WITH_DEVICE_IDVENDOR_INDEX => 0,
			STARTS_WITH_DEVICE_IDVENDOR_COUNT => 0,
			STARTS_WITH_DEVICE_IDPRODUCT_INDEX => 0,
			STARTS_WITH_DEVICE_IDPRODUCT_COUNT => 0,
			STARTS_WITH_DEVICE_BCDDEVICE_INDEX => 0,
			STARTS_WITH_DEVICE_BCDDEVICE_COUNT => 0,
			STARTS_WITH_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			STARTS_WITH_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			STARTS_WITH_DEVICE_IMANUFACTURER_INDEX => 0,
			STARTS_WITH_DEVICE_IMANUFACTURER_COUNT => 0,
			STARTS_WITH_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			STARTS_WITH_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			STARTS_WITH_DEVICE_IPRODUCT_INDEX => 0,
			STARTS_WITH_DEVICE_IPRODUCT_COUNT => 0,
			STARTS_WITH_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			STARTS_WITH_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			STARTS_WITH_DEVICE_ISERIALNUMBER_INDEX => 0,
			STARTS_WITH_DEVICE_ISERIALNUMBER_COUNT => 0,
			STARTS_WITH_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			STARTS_WITH_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			STARTS_WITH_CONFIGURATION_BLENGTH_INDEX => 0,
			STARTS_WITH_CONFIGURATION_BLENGTH_COUNT => 0,
			STARTS_WITH_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			STARTS_WITH_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			STARTS_WITH_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			STARTS_WITH_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			STARTS_WITH_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			STARTS_WITH_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			STARTS_WITH_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			STARTS_WITH_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			STARTS_WITH_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			STARTS_WITH_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			STARTS_WITH_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			STARTS_WITH_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			STARTS_WITH_CONFIGURATION_BMAXPOWER_INDEX => 0,
			STARTS_WITH_CONFIGURATION_BMAXPOWER_COUNT => 0,
			STARTS_WITH_INTERFACE_BLENGTH_INDEX => 0,
			STARTS_WITH_INTERFACE_BLENGTH_COUNT => 0,
			STARTS_WITH_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			STARTS_WITH_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			STARTS_WITH_INTERFACE_BALTERNATESETTING_INDEX => 0,
			STARTS_WITH_INTERFACE_BALTERNATESETTING_COUNT => 0,
			STARTS_WITH_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			STARTS_WITH_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			STARTS_WITH_INTERFACE_BINTERFACECLASS_INDEX => 0,
			STARTS_WITH_INTERFACE_BINTERFACECLASS_COUNT => 0,
			STARTS_WITH_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			STARTS_WITH_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			STARTS_WITH_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			STARTS_WITH_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			STARTS_WITH_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			STARTS_WITH_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			STARTS_WITH_INTERFACE_IINTERFACE_INDEX => 0,
			STARTS_WITH_INTERFACE_IINTERFACE_COUNT => 0,
			STARTS_WITH_HID_BLENGTH_INDEX => 0,
			STARTS_WITH_HID_BLENGTH_COUNT => 0,
			STARTS_WITH_HID_BCDHID_INDEX => 0,
			STARTS_WITH_HID_BCDHID_COUNT => 0,
			STARTS_WITH_HID_BCOUNTRYCODE_INDEX => 0,
			STARTS_WITH_HID_BCOUNTRYCODE_COUNT => 0,
			STARTS_WITH_HID_BNUMDESCRIPTORS_INDEX => 0,
			STARTS_WITH_HID_BNUMDESCRIPTORS_COUNT => 0,
			STARTS_WITH_HID_BDESCRIPTORTYPE_INDEX => 0,
			STARTS_WITH_HID_BDESCRIPTORTYPE_COUNT => 0,
			STARTS_WITH_HID_WDESCRIPTORLENGTH_INDEX => 0,
			STARTS_WITH_HID_WDESCRIPTORLENGTH_COUNT => 0,
			STARTS_WITH_ENDPOINT_BLENGTH_INDEX => 0,
			STARTS_WITH_ENDPOINT_BLENGTH_COUNT => 0,
			STARTS_WITH_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			STARTS_WITH_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			STARTS_WITH_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			STARTS_WITH_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			STARTS_WITH_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			STARTS_WITH_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			STARTS_WITH_ENDPOINT_BINTERVAL_INDEX => 0,
			STARTS_WITH_ENDPOINT_BINTERVAL_COUNT => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			STARTS_WITH_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			STARTS_WITH_OTHER_SPEED_BLENGTH_INDEX => 0,
			STARTS_WITH_OTHER_SPEED_BLENGTH_COUNT => 0,
			STARTS_WITH_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			STARTS_WITH_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			STARTS_WITH_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			STARTS_WITH_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			STARTS_WITH_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			STARTS_WITH_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			STARTS_WITH_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			STARTS_WITH_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			STARTS_WITH_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			STARTS_WITH_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			STARTS_WITH_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			STARTS_WITH_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			STARTS_WITH_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			STARTS_WITH_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			ENDS_WITH_MEMORY_ADDR_LENGTH => 1,
			ENDS_WITH_MEMORY_ADDR_MAX_INDEX => 0,
			ENDS_WITH_MEMORY_ADDR_MAX_COUNT => 0,
			ENDS_WITH_DEVICE_BLENGTH_INDEX => 0,
			ENDS_WITH_DEVICE_BLENGTH_COUNT => 0,
			ENDS_WITH_DEVICE_BCDUSB_INDEX => 0,
			ENDS_WITH_DEVICE_BCDUSB_COUNT => 0,
			ENDS_WITH_DEVICE_BDEVICECLASS_INDEX => 0,
			ENDS_WITH_DEVICE_BDEVICECLASS_COUNT => 0,
			ENDS_WITH_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			ENDS_WITH_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			ENDS_WITH_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			ENDS_WITH_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			ENDS_WITH_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			ENDS_WITH_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			ENDS_WITH_DEVICE_IDVENDOR_INDEX => 0,
			ENDS_WITH_DEVICE_IDVENDOR_COUNT => 0,
			ENDS_WITH_DEVICE_IDPRODUCT_INDEX => 0,
			ENDS_WITH_DEVICE_IDPRODUCT_COUNT => 0,
			ENDS_WITH_DEVICE_BCDDEVICE_INDEX => 0,
			ENDS_WITH_DEVICE_BCDDEVICE_COUNT => 0,
			ENDS_WITH_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			ENDS_WITH_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			ENDS_WITH_DEVICE_IMANUFACTURER_INDEX => 0,
			ENDS_WITH_DEVICE_IMANUFACTURER_COUNT => 0,
			ENDS_WITH_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			ENDS_WITH_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			ENDS_WITH_DEVICE_IPRODUCT_INDEX => 0,
			ENDS_WITH_DEVICE_IPRODUCT_COUNT => 0,
			ENDS_WITH_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			ENDS_WITH_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			ENDS_WITH_DEVICE_ISERIALNUMBER_INDEX => 0,
			ENDS_WITH_DEVICE_ISERIALNUMBER_COUNT => 0,
			ENDS_WITH_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			ENDS_WITH_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			ENDS_WITH_CONFIGURATION_BLENGTH_INDEX => 0,
			ENDS_WITH_CONFIGURATION_BLENGTH_COUNT => 0,
			ENDS_WITH_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			ENDS_WITH_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			ENDS_WITH_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			ENDS_WITH_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			ENDS_WITH_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			ENDS_WITH_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			ENDS_WITH_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			ENDS_WITH_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			ENDS_WITH_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			ENDS_WITH_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			ENDS_WITH_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			ENDS_WITH_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			ENDS_WITH_CONFIGURATION_BMAXPOWER_INDEX => 0,
			ENDS_WITH_CONFIGURATION_BMAXPOWER_COUNT => 0,
			ENDS_WITH_INTERFACE_BLENGTH_INDEX => 0,
			ENDS_WITH_INTERFACE_BLENGTH_COUNT => 0,
			ENDS_WITH_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			ENDS_WITH_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			ENDS_WITH_INTERFACE_BALTERNATESETTING_INDEX => 0,
			ENDS_WITH_INTERFACE_BALTERNATESETTING_COUNT => 0,
			ENDS_WITH_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			ENDS_WITH_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			ENDS_WITH_INTERFACE_BINTERFACECLASS_INDEX => 0,
			ENDS_WITH_INTERFACE_BINTERFACECLASS_COUNT => 0,
			ENDS_WITH_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			ENDS_WITH_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			ENDS_WITH_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			ENDS_WITH_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			ENDS_WITH_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			ENDS_WITH_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			ENDS_WITH_INTERFACE_IINTERFACE_INDEX => 0,
			ENDS_WITH_INTERFACE_IINTERFACE_COUNT => 0,
			ENDS_WITH_HID_BLENGTH_INDEX => 0,
			ENDS_WITH_HID_BLENGTH_COUNT => 0,
			ENDS_WITH_HID_BCDHID_INDEX => 0,
			ENDS_WITH_HID_BCDHID_COUNT => 0,
			ENDS_WITH_HID_BCOUNTRYCODE_INDEX => 0,
			ENDS_WITH_HID_BCOUNTRYCODE_COUNT => 0,
			ENDS_WITH_HID_BNUMDESCRIPTORS_INDEX => 0,
			ENDS_WITH_HID_BNUMDESCRIPTORS_COUNT => 0,
			ENDS_WITH_HID_BDESCRIPTORTYPE_INDEX => 0,
			ENDS_WITH_HID_BDESCRIPTORTYPE_COUNT => 0,
			ENDS_WITH_HID_WDESCRIPTORLENGTH_INDEX => 0,
			ENDS_WITH_HID_WDESCRIPTORLENGTH_COUNT => 0,
			ENDS_WITH_ENDPOINT_BLENGTH_INDEX => 0,
			ENDS_WITH_ENDPOINT_BLENGTH_COUNT => 0,
			ENDS_WITH_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			ENDS_WITH_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			ENDS_WITH_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			ENDS_WITH_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			ENDS_WITH_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			ENDS_WITH_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			ENDS_WITH_ENDPOINT_BINTERVAL_INDEX => 0,
			ENDS_WITH_ENDPOINT_BINTERVAL_COUNT => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			ENDS_WITH_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			ENDS_WITH_OTHER_SPEED_BLENGTH_INDEX => 0,
			ENDS_WITH_OTHER_SPEED_BLENGTH_COUNT => 0,
			ENDS_WITH_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			ENDS_WITH_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			ENDS_WITH_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			ENDS_WITH_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			ENDS_WITH_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			ENDS_WITH_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			ENDS_WITH_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			ENDS_WITH_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			ENDS_WITH_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			ENDS_WITH_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			ENDS_WITH_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			ENDS_WITH_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			ENDS_WITH_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			ENDS_WITH_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			CONTAINS_MEMORY_ADDR_LENGTH => 1,
			CONTAINS_MEMORY_ADDR_MAX_INDEX => 0,
			CONTAINS_MEMORY_ADDR_MAX_COUNT => 0,
			CONTAINS_DEVICE_BLENGTH_INDEX => 0,
			CONTAINS_DEVICE_BLENGTH_COUNT => 0,
			CONTAINS_DEVICE_BCDUSB_INDEX => 0,
			CONTAINS_DEVICE_BCDUSB_COUNT => 0,
			CONTAINS_DEVICE_BDEVICECLASS_INDEX => 0,
			CONTAINS_DEVICE_BDEVICECLASS_COUNT => 0,
			CONTAINS_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			CONTAINS_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			CONTAINS_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			CONTAINS_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			CONTAINS_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			CONTAINS_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			CONTAINS_DEVICE_IDVENDOR_INDEX => 0,
			CONTAINS_DEVICE_IDVENDOR_COUNT => 0,
			CONTAINS_DEVICE_IDPRODUCT_INDEX => 0,
			CONTAINS_DEVICE_IDPRODUCT_COUNT => 0,
			CONTAINS_DEVICE_BCDDEVICE_INDEX => 0,
			CONTAINS_DEVICE_BCDDEVICE_COUNT => 0,
			CONTAINS_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			CONTAINS_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			CONTAINS_DEVICE_IMANUFACTURER_INDEX => 0,
			CONTAINS_DEVICE_IMANUFACTURER_COUNT => 0,
			CONTAINS_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			CONTAINS_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			CONTAINS_DEVICE_IPRODUCT_INDEX => 0,
			CONTAINS_DEVICE_IPRODUCT_COUNT => 0,
			CONTAINS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			CONTAINS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			CONTAINS_DEVICE_ISERIALNUMBER_INDEX => 0,
			CONTAINS_DEVICE_ISERIALNUMBER_COUNT => 0,
			CONTAINS_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			CONTAINS_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			CONTAINS_CONFIGURATION_BLENGTH_INDEX => 0,
			CONTAINS_CONFIGURATION_BLENGTH_COUNT => 0,
			CONTAINS_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			CONTAINS_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			CONTAINS_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			CONTAINS_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			CONTAINS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			CONTAINS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			CONTAINS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			CONTAINS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			CONTAINS_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			CONTAINS_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			CONTAINS_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			CONTAINS_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			CONTAINS_CONFIGURATION_BMAXPOWER_INDEX => 0,
			CONTAINS_CONFIGURATION_BMAXPOWER_COUNT => 0,
			CONTAINS_INTERFACE_BLENGTH_INDEX => 0,
			CONTAINS_INTERFACE_BLENGTH_COUNT => 0,
			CONTAINS_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			CONTAINS_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			CONTAINS_INTERFACE_BALTERNATESETTING_INDEX => 0,
			CONTAINS_INTERFACE_BALTERNATESETTING_COUNT => 0,
			CONTAINS_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			CONTAINS_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			CONTAINS_INTERFACE_BINTERFACECLASS_INDEX => 0,
			CONTAINS_INTERFACE_BINTERFACECLASS_COUNT => 0,
			CONTAINS_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			CONTAINS_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			CONTAINS_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			CONTAINS_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			CONTAINS_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			CONTAINS_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			CONTAINS_INTERFACE_IINTERFACE_INDEX => 0,
			CONTAINS_INTERFACE_IINTERFACE_COUNT => 0,
			CONTAINS_HID_BLENGTH_INDEX => 0,
			CONTAINS_HID_BLENGTH_COUNT => 0,
			CONTAINS_HID_BCDHID_INDEX => 0,
			CONTAINS_HID_BCDHID_COUNT => 0,
			CONTAINS_HID_BCOUNTRYCODE_INDEX => 0,
			CONTAINS_HID_BCOUNTRYCODE_COUNT => 0,
			CONTAINS_HID_BNUMDESCRIPTORS_INDEX => 0,
			CONTAINS_HID_BNUMDESCRIPTORS_COUNT => 0,
			CONTAINS_HID_BDESCRIPTORTYPE_INDEX => 0,
			CONTAINS_HID_BDESCRIPTORTYPE_COUNT => 0,
			CONTAINS_HID_WDESCRIPTORLENGTH_INDEX => 0,
			CONTAINS_HID_WDESCRIPTORLENGTH_COUNT => 0,
			CONTAINS_ENDPOINT_BLENGTH_INDEX => 0,
			CONTAINS_ENDPOINT_BLENGTH_COUNT => 0,
			CONTAINS_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			CONTAINS_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			CONTAINS_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			CONTAINS_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			CONTAINS_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			CONTAINS_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			CONTAINS_ENDPOINT_BINTERVAL_INDEX => 0,
			CONTAINS_ENDPOINT_BINTERVAL_COUNT => 0,
			CONTAINS_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			CONTAINS_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			CONTAINS_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			CONTAINS_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			CONTAINS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			CONTAINS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			CONTAINS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			CONTAINS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			CONTAINS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			CONTAINS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			CONTAINS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			CONTAINS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			CONTAINS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			CONTAINS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			CONTAINS_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			CONTAINS_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			CONTAINS_OTHER_SPEED_BLENGTH_INDEX => 0,
			CONTAINS_OTHER_SPEED_BLENGTH_COUNT => 0,
			CONTAINS_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			CONTAINS_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			CONTAINS_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			CONTAINS_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			CONTAINS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			CONTAINS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			CONTAINS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			CONTAINS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			CONTAINS_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			CONTAINS_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			CONTAINS_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			CONTAINS_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			CONTAINS_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			CONTAINS_OTHER_SPEED_BMAXPOWER_COUNT => 0,

			NOT_CONTAINS_MEMORY_ADDR_LENGTH => 1,
			NOT_CONTAINS_MEMORY_ADDR_MAX_INDEX => 0,
			NOT_CONTAINS_MEMORY_ADDR_MAX_COUNT => 0,
			NOT_CONTAINS_DEVICE_BLENGTH_INDEX => 0,
			NOT_CONTAINS_DEVICE_BLENGTH_COUNT => 0,
			NOT_CONTAINS_DEVICE_BCDUSB_INDEX => 0,
			NOT_CONTAINS_DEVICE_BCDUSB_COUNT => 0,
			NOT_CONTAINS_DEVICE_BDEVICECLASS_INDEX => 0,
			NOT_CONTAINS_DEVICE_BDEVICECLASS_COUNT => 0,
			NOT_CONTAINS_DEVICE_BDEVICESUBCLASS_INDEX => 0,
			NOT_CONTAINS_DEVICE_BDEVICESUBCLASS_COUNT => 0,
			NOT_CONTAINS_DEVICE_BDEVICEPROTOCOL_INDEX => 0,
			NOT_CONTAINS_DEVICE_BDEVICEPROTOCOL_COUNT => 0,
			NOT_CONTAINS_DEVICE_BMAXPACKETSIZE0_INDEX => 0,
			NOT_CONTAINS_DEVICE_BMAXPACKETSIZE0_COUNT => 0,
			NOT_CONTAINS_DEVICE_IDVENDOR_INDEX => 0,
			NOT_CONTAINS_DEVICE_IDVENDOR_COUNT => 0,
			NOT_CONTAINS_DEVICE_IDPRODUCT_INDEX => 0,
			NOT_CONTAINS_DEVICE_IDPRODUCT_COUNT => 0,
			NOT_CONTAINS_DEVICE_BCDDEVICE_INDEX => 0,
			NOT_CONTAINS_DEVICE_BCDDEVICE_COUNT => 0,
			NOT_CONTAINS_DEVICE_IMANUFACTURER_BLENGTH_INDEX => 0,
			NOT_CONTAINS_DEVICE_IMANUFACTURER_BLENGTH_COUNT => 0,
			NOT_CONTAINS_DEVICE_IMANUFACTURER_INDEX => 0,
			NOT_CONTAINS_DEVICE_IMANUFACTURER_COUNT => 0,
			NOT_CONTAINS_DEVICE_IPRODUCT_BLENGTH_INDEX => 0,
			NOT_CONTAINS_DEVICE_IPRODUCT_BLENGTH_COUNT => 0,
			NOT_CONTAINS_DEVICE_IPRODUCT_INDEX => 0,
			NOT_CONTAINS_DEVICE_IPRODUCT_COUNT => 0,
			NOT_CONTAINS_DEVICE_ISERIALNUMBER_BLENGTH_INDEX => 0,
			NOT_CONTAINS_DEVICE_ISERIALNUMBER_BLENGTH_COUNT => 0,
			NOT_CONTAINS_DEVICE_ISERIALNUMBER_INDEX => 0,
			NOT_CONTAINS_DEVICE_ISERIALNUMBER_COUNT => 0,
			NOT_CONTAINS_DEVICE_BNUMCONFIGURATIONS_INDEX => 0,
			NOT_CONTAINS_DEVICE_BNUMCONFIGURATIONS_COUNT => 0,
			NOT_CONTAINS_CONFIGURATION_BLENGTH_INDEX => 0,
			NOT_CONTAINS_CONFIGURATION_BLENGTH_COUNT => 0,
			NOT_CONTAINS_CONFIGURATION_WTOTALLENGTH_INDEX => 0,
			NOT_CONTAINS_CONFIGURATION_WTOTALLENGTH_COUNT => 0,
			NOT_CONTAINS_CONFIGURATION_BNUMINTERFACES_INDEX => 0,
			NOT_CONTAINS_CONFIGURATION_BNUMINTERFACES_COUNT => 0,
			NOT_CONTAINS_CONFIGURATION_BCONFIGURATIONVALUE_INDEX => 0,
			NOT_CONTAINS_CONFIGURATION_BCONFIGURATIONVALUE_COUNT => 0,
			NOT_CONTAINS_CONFIGURATION_ICONFIGURATION_BLENGTH_INDEX => 0,
			NOT_CONTAINS_CONFIGURATION_ICONFIGURATION_BLENGTH_COUNT => 0,
			NOT_CONTAINS_CONFIGURATION_ICONFIGURATION_INDEX => 0,
			NOT_CONTAINS_CONFIGURATION_ICONFIGURATION_COUNT => 0,
			NOT_CONTAINS_CONFIGURATION_BMATTRIBUTES_INDEX => 0,
			NOT_CONTAINS_CONFIGURATION_BMATTRIBUTES_COUNT => 0,
			NOT_CONTAINS_CONFIGURATION_BMAXPOWER_INDEX => 0,
			NOT_CONTAINS_CONFIGURATION_BMAXPOWER_COUNT => 0,
			NOT_CONTAINS_INTERFACE_BLENGTH_INDEX => 0,
			NOT_CONTAINS_INTERFACE_BLENGTH_COUNT => 0,
			NOT_CONTAINS_INTERFACE_BINTERFACENUMBER_INDEX => 0,
			NOT_CONTAINS_INTERFACE_BINTERFACENUMBER_COUNT => 0,
			NOT_CONTAINS_INTERFACE_BALTERNATESETTING_INDEX => 0,
			NOT_CONTAINS_INTERFACE_BALTERNATESETTING_COUNT => 0,
			NOT_CONTAINS_INTERFACE_BNUMENDPOINTS_INDEX => 0,
			NOT_CONTAINS_INTERFACE_BNUMENDPOINTS_COUNT => 0,
			NOT_CONTAINS_INTERFACE_BINTERFACECLASS_INDEX => 0,
			NOT_CONTAINS_INTERFACE_BINTERFACECLASS_COUNT => 0,
			NOT_CONTAINS_INTERFACE_BINTERFACESUBCLASS_INDEX => 0,
			NOT_CONTAINS_INTERFACE_BINTERFACESUBCLASS_COUNT => 0,
			NOT_CONTAINS_INTERFACE_BINTERFACEPROTOCOL_INDEX => 0,
			NOT_CONTAINS_INTERFACE_BINTERFACEPROTOCOL_COUNT => 0,
			NOT_CONTAINS_INTERFACE_IINTERFACE_BLENGTH_INDEX => 0,
			NOT_CONTAINS_INTERFACE_IINTERFACE_BLENGTH_COUNT => 0,
			NOT_CONTAINS_INTERFACE_IINTERFACE_INDEX => 0,
			NOT_CONTAINS_INTERFACE_IINTERFACE_COUNT => 0,
			NOT_CONTAINS_HID_BLENGTH_INDEX => 0,
			NOT_CONTAINS_HID_BLENGTH_COUNT => 0,
			NOT_CONTAINS_HID_BCDHID_INDEX => 0,
			NOT_CONTAINS_HID_BCDHID_COUNT => 0,
			NOT_CONTAINS_HID_BCOUNTRYCODE_INDEX => 0,
			NOT_CONTAINS_HID_BCOUNTRYCODE_COUNT => 0,
			NOT_CONTAINS_HID_BNUMDESCRIPTORS_INDEX => 0,
			NOT_CONTAINS_HID_BNUMDESCRIPTORS_COUNT => 0,
			NOT_CONTAINS_HID_BDESCRIPTORTYPE_INDEX => 0,
			NOT_CONTAINS_HID_BDESCRIPTORTYPE_COUNT => 0,
			NOT_CONTAINS_HID_WDESCRIPTORLENGTH_INDEX => 0,
			NOT_CONTAINS_HID_WDESCRIPTORLENGTH_COUNT => 0,
			NOT_CONTAINS_ENDPOINT_BLENGTH_INDEX => 0,
			NOT_CONTAINS_ENDPOINT_BLENGTH_COUNT => 0,
			NOT_CONTAINS_ENDPOINT_BENDPOINTADDRESS_INDEX => 0,
			NOT_CONTAINS_ENDPOINT_BENDPOINTADDRESS_COUNT => 0,
			NOT_CONTAINS_ENDPOINT_BMATTRIBUTES_INDEX => 0,
			NOT_CONTAINS_ENDPOINT_BMATTRIBUTES_COUNT => 0,
			NOT_CONTAINS_ENDPOINT_WMAXPACKETSIZE_INDEX => 0,
			NOT_CONTAINS_ENDPOINT_WMAXPACKETSIZE_COUNT => 0,
			NOT_CONTAINS_ENDPOINT_BINTERVAL_INDEX => 0,
			NOT_CONTAINS_ENDPOINT_BINTERVAL_COUNT => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BLENGTH_INDEX => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BLENGTH_COUNT => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BCDUSB_INDEX => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BCDUSB_COUNT => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICECLASS_INDEX => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICECLASS_COUNT => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICESUBCLASS_INDEX => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICESUBCLASS_COUNT => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_INDEX => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BDEVICEPROTOCOL_COUNT => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_INDEX => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BMAXPACKETSIZE0_COUNT => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_INDEX => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BNUMCONFIGURATIONS_COUNT => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BRESERVED_INDEX => 0,
			NOT_CONTAINS_DEVICE_QUALIFIER_BRESERVED_COUNT => 0,
			NOT_CONTAINS_OTHER_SPEED_BLENGTH_INDEX => 0,
			NOT_CONTAINS_OTHER_SPEED_BLENGTH_COUNT => 0,
			NOT_CONTAINS_OTHER_SPEED_WTOTALLENGTH_INDEX => 0,
			NOT_CONTAINS_OTHER_SPEED_WTOTALLENGTH_COUNT => 0,
			NOT_CONTAINS_OTHER_SPEED_BNUMINTERFACES_INDEX => 0,
			NOT_CONTAINS_OTHER_SPEED_BNUMINTERFACES_COUNT => 0,
			NOT_CONTAINS_OTHER_SPEED_BCONFIGURATIONVALUE_INDEX => 0,
			NOT_CONTAINS_OTHER_SPEED_BCONFIGURATIONVALUE_COUNT => 0,
			NOT_CONTAINS_OTHER_SPEED_ICONFIGURATION_BLENGTH_INDEX => 0,
			NOT_CONTAINS_OTHER_SPEED_ICONFIGURATION_BLENGTH_COUNT => 0,
			NOT_CONTAINS_OTHER_SPEED_ICONFIGURATION_INDEX => 0,
			NOT_CONTAINS_OTHER_SPEED_ICONFIGURATION_COUNT => 0,
			NOT_CONTAINS_OTHER_SPEED_BMATTRIBUTES_INDEX => 0,
			NOT_CONTAINS_OTHER_SPEED_BMATTRIBUTES_COUNT => 0,
			NOT_CONTAINS_OTHER_SPEED_BMAXPOWER_INDEX => 0,
			NOT_CONTAINS_OTHER_SPEED_BMAXPOWER_COUNT => 0
		)

		PORT MAP (
			i_sys_clock => i_sys_clock,
			i_enable => i_enable,
			i_descriptor_field => i_descriptor_field,
			i_descriptor_field_available => i_descriptor_field_available,
			i_descriptor_value => i_descriptor_value,
			i_descriptor_value_en => i_descriptor_value_en,
			i_descriptor_value_total_part_number => i_descriptor_value_total_part_number,
			i_descriptor_value_part_number => i_descriptor_value_part_number,
			i_descriptor_value_new_part => i_descriptor_value_new_part,
			o_descriptor_value_next_part_request => o_descriptor_value_next_part_request,
			o_ready => o_ready,
			o_result => o_result
	);

end Behavioral;
