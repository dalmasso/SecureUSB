------------------------------------------------------------------------
-- Engineer:    Dalmasso Loic
-- Create Date: 30/07/2025
-- Package Name: USBDescriptorFields
-- Description:
--		Package assigning USB Descriptor Fields to unique values
------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE USBDescriptorFields is

	-- USB Descriptor Field Length
	constant USB_DESCRIPTOR_FIELD_BIT_LENGTH: INTEGER := 12;

	-- Device Descriptor (0x01)
	constant DEVICE_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"010";
	constant DEVICE_BCDUSB_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"011";
	constant DEVICE_BDEVICECLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"012";
	constant DEVICE_BDEVICESUBCLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"013";
	constant DEVICE_BDEVICEPROTOCOL_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"014";
	constant DEVICE_BMAXPACKETSIZE0_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"015";
	constant DEVICE_IDVENDOR_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"016";
	constant DEVICE_IDPRODUCT_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"017";
	constant DEVICE_BCDDEVICE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"018";
	constant DEVICE_BNUMCONFIGURATIONS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"019";

	-- Device Qualifier Descriptor (0x06)
	constant DEVICE_QUALIFIER_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"060";
	constant DEVICE_QUALIFIER_BCDUSB_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"061";
	constant DEVICE_QUALIFIER_BDEVICECLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"062";
	constant DEVICE_QUALIFIER_BDEVICESUBCLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"063";
	constant DEVICE_QUALIFIER_BDEVICEPROTOCOL_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"064";
	constant DEVICE_QUALIFIER_BMAXPACKETSIZE0_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"065";
	constant DEVICE_QUALIFIER_BCDDEVICE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"066";
	constant DEVICE_QUALIFIER_BNUMCONFIGURATIONS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"067";
	constant DEVICE_QUALIFIER_BRESERVED_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"068";

	-- Configuration Descriptor (0x02)
	constant CONFIGURATION_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"020";
	constant CONFIGURATION_WTOTALLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"021";
	constant CONFIGURATION_BNUMINTERFACES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"022";
	constant CONFIGURATION_BCONFIGURATIONVALUE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"023";
	constant CONFIGURATION_BMATTRIBUTES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"024";
	constant CONFIGURATION_BMAXPOWER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"025";

	-- Other Speed Descriptor (0x07)
	constant OTHER_SPEED_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"070";
	constant OTHER_SPEED_WTOTALLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"071";
	constant OTHER_SPEED_BNUMINTERFACES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"072";
	constant OTHER_SPEED_BCONFIGURATIONVALUE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"073";
	constant OTHER_SPEED_BMATTRIBUTES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"074";
	constant OTHER_SPEED_BMAXPOWER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"075";

	-- Interface Descriptor (0x04)
	constant INTERFACE_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"040";
	constant INTERFACE_BINTERFACENUMBER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"041";
	constant INTERFACE_BALTERNATESETTING_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"042";
	constant INTERFACE_BNUMENDPOINTS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"043";
	constant INTERFACE_BINTERFACECLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"044";
	constant INTERFACE_BINTERFACESUBCLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"045";
	constant INTERFACE_BINTERFACEPROTOCOL_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"046";

	-- Endpoint Descriptor (0x05)
	constant ENDPOINT_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"050";
	constant ENDPOINT_BENDPOINTADDRESS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"051";
	constant ENDPOINT_BMATTRIBUTES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"052";
	constant ENDPOINT_WMAXPACKETSIZE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"053";
	constant ENDPOINT_BINTERVAL_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"054";

	-- HID Descriptor (0x21)
	constant HID_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"210";
	constant HID_BCDHID_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"211";
	constant HID_BCOUNTRYCODE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"212";
	constant HID_BNUMDESCRIPTORS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"213";
	constant HID_BDESCRIPTORTYPE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"214";
	constant HID_WDESCRIPTORLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"215";

	-- String Descriptor (0x03)
	constant STRING_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"030";
	constant STRING_IMANUFACTURER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"031";
	constant STRING_IPRODUCT_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"032";
	constant STRING_ISERIALNUMBER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"033";
	constant STRING_ICONFIGURATION_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"034";
	constant STRING_IINTERFACE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"035";

END PACKAGE USBDescriptorFields;