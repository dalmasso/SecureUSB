------------------------------------------------------------------------
-- Engineer:    Dalmasso Loic
-- Create Date: 30/07/2025
-- Package Name: USBDescriptorFields
-- Description:
--		Package assigning USB Descriptor Fields to unique values
------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE USBDescriptorFields is

	-- USB Descriptor Field Length
	constant USB_DESCRIPTOR_FIELD_BIT_LENGTH: INTEGER := 12;

	-- USB Descriptor Request Types
	constant USB_DESCRIPTOR_DEVICE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"001";
	constant USB_DESCRIPTOR_CONFIGURATION_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"002";
	constant USB_DESCRIPTOR_STRING_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"003";
	constant USB_DESCRIPTOR_INTERFACE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"004";
	constant USB_DESCRIPTOR_ENDPOINT_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"005";
	constant USB_DESCRIPTOR_DEVICE_QUALIFIER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"006";
	constant USB_DESCRIPTOR_OTHER_SPEED_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"007";
	constant USB_DESCRIPTOR_HID_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"021";

	-- Device Descriptor (0x01)
	constant DEVICE_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"010";
	constant DEVICE_BCDUSB_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"011";
	constant DEVICE_BDEVICECLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"012";
	constant DEVICE_BDEVICESUBCLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"013";
	constant DEVICE_BDEVICEPROTOCOL_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"014";
	constant DEVICE_BMAXPACKETSIZE0_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"015";
	constant DEVICE_IDVENDOR_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"016";
	constant DEVICE_IDPRODUCT_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"017";
	constant DEVICE_BCDDEVICE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"018";
	constant DEVICE_IMANUFACTURER_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"019";
	constant DEVICE_IMANUFACTURER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"01A";
	constant DEVICE_IPRODUCT_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"01B";
	constant DEVICE_IPRODUCT_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"01C";
	constant DEVICE_ISERIALNUMBER_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"01D";
	constant DEVICE_ISERIALNUMBER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"01E";
	constant DEVICE_BNUMCONFIGURATIONS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"01F";

	-- Configuration Descriptor (0x02)
	constant CONFIGURATION_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"020";
	constant CONFIGURATION_WTOTALLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"021";
	constant CONFIGURATION_BNUMINTERFACES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"022";
	constant CONFIGURATION_BCONFIGURATIONVALUE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"023";
	constant CONFIGURATION_ICONFIGURATION_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"024";
	constant CONFIGURATION_ICONFIGURATION_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"025";	
	constant CONFIGURATION_BMATTRIBUTES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"026";
	constant CONFIGURATION_BMAXPOWER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"027";

	-- Interface Descriptor (0x04)
	constant INTERFACE_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"040";
	constant INTERFACE_BINTERFACENUMBER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"041";
	constant INTERFACE_BALTERNATESETTING_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"042";
	constant INTERFACE_BNUMENDPOINTS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"043";
	constant INTERFACE_BINTERFACECLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"044";
	constant INTERFACE_BINTERFACESUBCLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"045";
	constant INTERFACE_BINTERFACEPROTOCOL_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"046";
	constant INTERFACE_IINTERFACE_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"047";
	constant INTERFACE_IINTERFACE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"048";

    -- HID Descriptor (0x21)
	constant HID_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"210";
	constant HID_BCDHID_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"211";
	constant HID_BCOUNTRYCODE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"212";
	constant HID_BNUMDESCRIPTORS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"213";
	constant HID_BDESCRIPTORTYPE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"214";
	constant HID_WDESCRIPTORLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"215";

	-- Endpoint Descriptor (0x05)
	constant ENDPOINT_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"050";
	constant ENDPOINT_BENDPOINTADDRESS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"051";
	constant ENDPOINT_BMATTRIBUTES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"052";
	constant ENDPOINT_WMAXPACKETSIZE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"053";
	constant ENDPOINT_BINTERVAL_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"054";

    -- Device Qualifier Descriptor (0x06)
	constant DEVICE_QUALIFIER_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"060";
	constant DEVICE_QUALIFIER_BCDUSB_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"061";
	constant DEVICE_QUALIFIER_BDEVICECLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"062";
	constant DEVICE_QUALIFIER_BDEVICESUBCLASS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"063";
	constant DEVICE_QUALIFIER_BDEVICEPROTOCOL_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"064";
	constant DEVICE_QUALIFIER_BMAXPACKETSIZE0_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"065";
	constant DEVICE_QUALIFIER_BCDDEVICE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"066";
	constant DEVICE_QUALIFIER_BNUMCONFIGURATIONS_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"067";
	constant DEVICE_QUALIFIER_BRESERVED_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"068";

	-- Other Speed Descriptor (0x07)
	constant OTHER_SPEED_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"070";
	constant OTHER_SPEED_WTOTALLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"071";
	constant OTHER_SPEED_BNUMINTERFACES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"072";
	constant OTHER_SPEED_BCONFIGURATIONVALUE_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"073";
	constant OTHER_SPEED_ICONFIGURATION_BLENGTH_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"074";
	constant OTHER_SPEED_ICONFIGURATION_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"075";	
	constant OTHER_SPEED_BMATTRIBUTES_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"076";
	constant OTHER_SPEED_BMAXPOWER_TYPE: UNSIGNED(USB_DESCRIPTOR_FIELD_BIT_LENGTH-1 downto 0) := x"077";

END PACKAGE USBDescriptorFields;
